`include "..\src\Top_example.sv"
//`include "Random.sv"
`include "..\src\DE2_115/SevenHexDecoder.sv"
`include "..\src\DE2_115/Debounce.sv"
`include "..\src\DE2_115/DE2_115.sv"
